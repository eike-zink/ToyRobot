module main

import toy_robot

fn main() {
	robot := toy_robot.Robot{ name: 'Tobi' }

	println('Hello $robot.name')

}
